
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--use IEEE.STD_LOGIC_ARITH.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity display is
    Port(  
        ins_value, wd_out: in std_logic_vector(31 downto 0);
        mode: in std_logic_vector(3 downto 0);
        pc, rf_value: in std_logic_vector(31 downto 0);
        led1,led2,led3,led4,led5,led6,led7,led8,led9,led10,led11,led12,led13,led14,led15,led16:out std_logic;
        state_out: in std_logic_vector(6 downto 0);
        IR_in, DR_in, A_in, B_in, RES_in: in std_logic_vector(31 downto 0);
        z_in, c_in, v_in, n_in: in std_logic
    );
end display;

architecture Behavioral of display is
begin
	process(mode, wd_out, ins_value, IR_in, DR_in, A_in, B_in, RES_in, pc, rf_value, state_out, z_in, n_in, c_in, v_in)
	begin
        led1<='0';
        led2<='0';
        led3<='0';
        led4<='0';
        led5<='0';
        led6<='0';
        led7<='0';
        led8<='0';
        led9<='0';
        led10<='0';
        led11<='0';
        led12<='0';
        led13<='0';
        led14<='0';
        led15<='0';
        led16 <= '0';
		case mode is
			when "0000"=> -- Data written to the DM
--				if (wd_out(0)='1') then led1<='1'; end if;
--				if (wd_out(1)='1') then led2<='1'; end if;
--				if (wd_out(2)='1') then led3<='1'; end if;
--				if (wd_out(3)='1') then led4<='1'; end if;
--				if (wd_out(4)='1') then led5<='1'; end if;
--				if (wd_out(5)='1') then led6<='1'; end if;
--				if (wd_out(6)='1') then led7<='1'; end if;
--				if (wd_out(7)='1') then led8<='1'; end if;
--				if (wd_out(8)='1') then led9<='1'; end if;
--				if (wd_out(9)='1') then led10<='1'; end if;
--				if (wd_out(10)='1') then led11<='1'; end if;
--				if (wd_out(11)='1') then led12<='1'; end if;
--				if (wd_out(12)='1') then led13<='1'; end if;
--				if (wd_out(13)='1') then led14<='1'; end if;
--				if (wd_out(14)='1') then led15<='1'; end if;
--				if (wd_out(15)='1') then led16<='1'; end if;
                if IR_in(16) = '1' then led1 <= '1'; end if;
                if IR_in(17) = '1' then led2 <= '1'; end if;
                if IR_in(18) = '1' then led3 <= '1'; end if;
                if IR_in(19) = '1' then led4 <= '1'; end if;
                if IR_in(20) = '1' then led5 <= '1'; end if;
                if IR_in(21) = '1' then led6 <= '1'; end if;
                if IR_in(22) = '1' then led7 <= '1'; end if;
                if IR_in(23) = '1' then led8 <= '1'; end if;
                if IR_in(24) = '1' then led9 <= '1'; end if;
                if IR_in(25) = '1' then led10 <= '1'; end if;
                if IR_in(26) = '1' then led11 <= '1'; end if;
                if IR_in(27) = '1' then led12 <= '1'; end if;
                if IR_in(28) = '1' then led13 <= '1'; end if;
                if IR_in(29) = '1' then led14 <= '1'; end if;
                if IR_in(30) = '1' then led15 <= '1'; end if;
                if IR_in(31) = '1' then led16 <= '1'; end if;
			when "0001"=> -- Value of Rn
--				if (ins_value(16)='1') then led1<='1';end if;
--				if (ins_value(17)='1') then led2<='1';end if;
--				if (ins_value(18)='1') then led3<='1';end if;
--				if (ins_value(19)='1') then led4<='1';end if;
                if A_in(0) = '1' then led1 <= '1'; end if;
                if A_in(1) = '1' then led2 <= '1'; end if;
                if A_in(2) = '1' then led3 <= '1'; end if;
                if A_in(3) = '1' then led4 <= '1'; end if;
                if A_in(4) = '1' then led5 <= '1'; end if;
                if A_in(5) = '1' then led6 <= '1'; end if;
                if A_in(6) = '1' then led7 <= '1'; end if;
                if A_in(7) = '1' then led8 <= '1'; end if;
                if A_in(8) = '1' then led9 <= '1'; end if;
                if A_in(9) = '1' then led10 <= '1'; end if;
                if A_in(10) = '1' then led11 <= '1'; end if;
                if A_in(11) = '1' then led12 <= '1'; end if;
                if A_in(12) = '1' then led13 <= '1'; end if;
                if A_in(13) = '1' then led14 <= '1'; end if;
                if A_in(14) = '1' then led15 <= '1'; end if;
                if A_in(15) = '1' then led16 <= '1'; end if;
			when "0010"=> -- Value of Rd
--				if (ins_value(15)='1') then led1<='1';end if;
--				if (ins_value(14)='1') then led2<='1';end if;
--				if (ins_value(13)='1') then led3<='1';end if;
--				if (ins_value(12)='1') then led4<='1';end if;
                if B_in(0) = '1' then led1 <= '1'; end if;
                if B_in(1) = '1' then led2 <= '1'; end if;
                if B_in(2) = '1' then led3 <= '1'; end if;
                if B_in(3) = '1' then led4 <= '1'; end if;
                if B_in(4) = '1' then led5 <= '1'; end if;
                if B_in(5) = '1' then led6 <= '1'; end if;
                if B_in(6) = '1' then led7 <= '1'; end if;
                if B_in(7) = '1' then led8 <= '1'; end if;
                if B_in(8) = '1' then led9 <= '1'; end if;
                if B_in(9) = '1' then led10 <= '1'; end if;
                if B_in(10) = '1' then led11 <= '1'; end if;
                if B_in(11) = '1' then led12 <= '1'; end if;
                if B_in(12) = '1' then led13 <= '1'; end if;
                if B_in(13) = '1' then led14 <= '1'; end if;
                if B_in(14) = '1' then led15 <= '1'; end if;
                if B_in(15) = '1' then led16 <= '1'; end if;
			when "0011"=> -- Cond
--				if (ins_value(28)='1') then led1<='1';end if;
--				if (ins_value(29)='1') then led2<='1';end if;
--				if (ins_value(30)='1') then led3<='1';end if;
--				if (ins_value(31)='1') then led4<='1';end if;
                if RES_in(0) = '1' then led1 <= '1'; end if;
                if RES_in(1) = '1' then led2 <= '1'; end if;
                if RES_in(2) = '1' then led3 <= '1'; end if;
                if RES_in(3) = '1' then led4 <= '1'; end if;
                if RES_in(4) = '1' then led5 <= '1'; end if;
                if RES_in(5) = '1' then led6 <= '1'; end if;
                if RES_in(6) = '1' then led7 <= '1'; end if;
                if RES_in(7) = '1' then led8 <= '1'; end if;
                if RES_in(8) = '1' then led9 <= '1'; end if;
                if RES_in(9) = '1' then led10 <= '1'; end if;
                if RES_in(10) = '1' then led11 <= '1'; end if;
                if RES_in(11) = '1' then led12 <= '1'; end if;
                if RES_in(12) = '1' then led13 <= '1'; end if;
                if RES_in(13) = '1' then led14 <= '1'; end if;
                if RES_in(14) = '1' then led15 <= '1'; end if;
                if RES_in(15) = '1' then led16 <= '1'; end if;
			when "0100"=> -- Second operand
--				if (ins_value(0)='1') then led1<='1'; end if;
--				if (ins_value(1)='1') then led2<='1'; end if;
--				if (ins_value(2)='1') then led3<='1'; end if;
--				if (ins_value(3)='1') then led4<='1'; end if;
--				if (ins_value(4)='1') then led5<='1'; end if;
--				if (ins_value(5)='1') then led6<='1'; end if;
--				if (ins_value(6)='1') then led7<='1'; end if;
--				if (ins_value(7)='1') then led8<='1'; end if;
--				if (ins_value(8)='1') then led9<='1'; end if;
--				if (ins_value(9)='1') then led10<='1'; end if;
--				if (ins_value(10)='1') then led11<='1'; end if;
--				if (ins_value(11)='1') then led12<='1'; end if;
                if DR_in(0) = '1' then led1 <= '1'; end if;
                if DR_in(1) = '1' then led2 <= '1'; end if;
                if DR_in(2) = '1' then led3 <= '1'; end if;
                if DR_in(3) = '1' then led4 <= '1'; end if;
                if DR_in(4) = '1' then led5 <= '1'; end if;
                if DR_in(5) = '1' then led6 <= '1'; end if;
                if DR_in(6) = '1' then led7 <= '1'; end if;
                if DR_in(7) = '1' then led8 <= '1'; end if;
                if DR_in(8) = '1' then led9 <= '1'; end if;
                if DR_in(9) = '1' then led10 <= '1'; end if;
                if DR_in(10) = '1' then led11 <= '1'; end if;
                if DR_in(11) = '1' then led12 <= '1'; end if;
                if DR_in(12) = '1' then led13 <= '1'; end if;
                if DR_in(13) = '1' then led14 <= '1'; end if;
                if DR_in(14) = '1' then led15 <= '1'; end if;
                if DR_in(15) = '1' then led16 <= '1'; end if;
            when "1000" => -- Lower 16 bits of ins_value
                led1 <= ins_value(0);
                led2 <= ins_value(1);
                led3 <= ins_value(2);
                led4 <= ins_value(3);
                led5 <= ins_value(4);
                led6 <= ins_value(5);
                led7 <= ins_value(6);
                led8 <= ins_value(7);
                led9 <= ins_value(8);
                led10 <= ins_value(9);
                led11 <= ins_value(10);
                led12 <= ins_value(11);
                led13 <= ins_value(12);
                led14 <= ins_value(13);
                led15 <= ins_value(14);
                led16 <= ins_value(15);
            when "1001" =>
                led1 <= ins_value(16);
                led2 <= ins_value(17);
                led3 <= ins_value(18);
                led4 <= ins_value(19);
                led5 <= ins_value(20);
                led6 <= ins_value(21);
                led7 <= ins_value(22);
                led8 <= ins_value(23);
                led9 <= ins_value(24);
                led10 <= ins_value(25);
                led11 <= ins_value(26);
                led12 <= ins_value(27);
                led13 <= ins_value(28);
                led14 <= ins_value(29);
                led15 <= ins_value(30);
                led16 <= ins_value(31);
            when "1010" =>
                led1 <= pc(0);
                led2 <= pc(1);
                led3 <= pc(2);
                led4 <= pc(3);
                led5 <= pc(4);
                led6 <= pc(5);
                led7 <= pc(6);
                led8 <= pc(7);
                led9 <= pc(8);
                led10 <= pc(9);
                led11 <= pc(10);
                led12 <= pc(11);
                led13 <= pc(12);
                led14 <= pc(13);
                led15 <= pc(14);
                led16 <= pc(15);
            when "1011" =>
                led1 <= rf_value(0);
                led2 <= rf_value(1);
                led3 <= rf_value(2);
                led4 <= rf_value(3);
                led5 <= rf_value(4);
                led6 <= rf_value(5);
                led7 <= rf_value(6);
                led8 <= rf_value(7);
                led9 <= rf_value(8);
                led10 <= rf_value(9);
                led11 <= rf_value(10);
                led12 <= rf_value(11);
                led13 <= rf_value(12);
                led14 <= rf_value(13);
                led15 <= rf_value(14);
                led16 <= rf_value(15);
            when "1100" =>
                led1 <= state_out(0);
                led2 <= state_out(1);
                led3 <= state_out(2);
                led4 <= state_out(3);
                led5<= z_in;
                led6<= n_in;
                led7<= c_in;
                led8<= v_in;
                led9<='0';
                led10<='0';
                led11<='0';
                led12<='0';
                led13<='0';
                led14<=state_out(4);
                led15<=state_out(5);
                led16 <= state_out(6);
         when others=>
                led1<='0';
                led2<='0';
                led3<='0';
                led4<='0';
                led5<='0';
                led6<='0';
                led7<='0';
                led8<='0';
                led9<='0';
                led10<='0';
                led11<='0';
                led12<='0';
                led13<='0';
                led14<='0';
                led15<='0';
                led16 <= '0';
		end case;
	end process;
end architecture;
